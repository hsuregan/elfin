module crc8_byte_tb;
